`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:46:28 05/16/2022 
// Design Name: 
// Module Name:    C1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module C1(eqz1,neqz1,z);
input z;
output reg eqz,neqz;
always@(posedge clk)
if(z) ==0;


endmodule
